// SuperRT by Ben Carter (c) 2021
// Character data ROM for debug display

`include "Config.sv"

module CharROM (
	input [3:0] char,
	input [2:0] x,
	input [2:0] y,
	
	output [0:0] pixel
);

// Bitmaps
reg [7:0] data[128];

assign pixel = (data[{ char, y }] >> (7 - x));

initial begin
	data[  0] = 8'b00000000;
	data[  1] = 8'b00000000;
	data[  2] = 8'b01111110;
	data[  3] = 8'b01000010;
	data[  4] = 8'b01000010;
	data[  5] = 8'b01000010;
	data[  6] = 8'b01111110;
	data[  7] = 8'b00000000;
	
	data[  8] = 8'b00000000;
	data[  9] = 8'b00000000;
	data[ 10] = 8'b00010000;
	data[ 11] = 8'b00010000;
	data[ 12] = 8'b00010000;
	data[ 13] = 8'b00010000;
	data[ 14] = 8'b00010000;
	data[ 15] = 8'b00000000;

	data[ 16] = 8'b00000000;
	data[ 17] = 8'b00000000;
	data[ 18] = 8'b01111110;
	data[ 19] = 8'b00000010;
	data[ 20] = 8'b01111110;
	data[ 21] = 8'b01000000;
	data[ 22] = 8'b01111110;
	data[ 23] = 8'b00000000;

	data[ 24] = 8'b00000000;
	data[ 25] = 8'b00000000;
	data[ 26] = 8'b01111110;
	data[ 27] = 8'b00000010;
	data[ 28] = 8'b00011110;
	data[ 29] = 8'b00000010;
	data[ 30] = 8'b01111110;
	data[ 31] = 8'b00000000;

	data[ 32] = 8'b00000000;
	data[ 33] = 8'b00000000;
	data[ 34] = 8'b01001000;
	data[ 35] = 8'b01001000;
	data[ 36] = 8'b01001000;
	data[ 37] = 8'b01111110;
	data[ 38] = 8'b00001000;
	data[ 39] = 8'b00000000;

	data[ 40] = 8'b00000000;
	data[ 41] = 8'b00000000;
	data[ 42] = 8'b01111110;
	data[ 43] = 8'b01000000;
	data[ 44] = 8'b01111110;
	data[ 45] = 8'b00000010;
	data[ 46] = 8'b01111110;
	data[ 47] = 8'b00000000;

	data[ 48] = 8'b00000000;
	data[ 49] = 8'b00000000;
	data[ 50] = 8'b01000000;
	data[ 51] = 8'b01000000;
	data[ 52] = 8'b01111110;
	data[ 53] = 8'b01000010;
	data[ 54] = 8'b01111110;
	data[ 55] = 8'b00000000;

	data[ 56] = 8'b00000000;
	data[ 57] = 8'b00000000;
	data[ 58] = 8'b00111110;
	data[ 59] = 8'b00000010;
	data[ 60] = 8'b00000010;
	data[ 61] = 8'b00000010;
	data[ 62] = 8'b00000010;
	data[ 63] = 8'b00000000;

	data[ 64] = 8'b00000000;
	data[ 65] = 8'b00000000;
	data[ 66] = 8'b01111110;
	data[ 67] = 8'b01000010;
	data[ 68] = 8'b01111110;
	data[ 69] = 8'b01000010;
	data[ 70] = 8'b01111110;
	data[ 71] = 8'b00000000;

	data[ 72] = 8'b00000000;
	data[ 73] = 8'b00000000;
	data[ 74] = 8'b01111110;
	data[ 75] = 8'b01000010;
	data[ 76] = 8'b01111110;
	data[ 77] = 8'b00000010;
	data[ 78] = 8'b01111110;
	data[ 79] = 8'b00000000;

	data[ 80] = 8'b00000000;
	data[ 81] = 8'b00000000;
	data[ 82] = 8'b00111100;
	data[ 83] = 8'b01000010;
	data[ 84] = 8'b01111110;
	data[ 85] = 8'b01000010;
	data[ 86] = 8'b01000010;
	data[ 87] = 8'b00000000;

	data[ 88] = 8'b00000000;
	data[ 89] = 8'b00000000;
	data[ 90] = 8'b01111100;
	data[ 91] = 8'b01000010;
	data[ 92] = 8'b01111100;
	data[ 93] = 8'b01000010;
	data[ 94] = 8'b01111100;
	data[ 95] = 8'b00000000;

	data[ 96] = 8'b00000000;
	data[ 97] = 8'b00000000;
	data[ 98] = 8'b01111110;
	data[ 99] = 8'b01000000;
	data[100] = 8'b01000000;
	data[101] = 8'b01000000;
	data[102] = 8'b01111110;
	data[103] = 8'b00000000;

	data[104] = 8'b00000000;
	data[105] = 8'b00000000;
	data[106] = 8'b01111100;
	data[107] = 8'b01000010;
	data[108] = 8'b01000010;
	data[109] = 8'b01000010;
	data[110] = 8'b01111100;
	data[111] = 8'b00000000;

	data[112] = 8'b00000000;
	data[113] = 8'b00000000;
	data[114] = 8'b01111110;
	data[115] = 8'b01000000;
	data[116] = 8'b01110000;
	data[117] = 8'b01000000;
	data[118] = 8'b01111110;
	data[119] = 8'b00000000;

	data[120] = 8'b00000000;
	data[121] = 8'b00000000;
	data[122] = 8'b01111110;
	data[123] = 8'b01000000;
	data[124] = 8'b01111110;
	data[125] = 8'b01000000;
	data[126] = 8'b01000000;
	data[127] = 8'b00000000;
end

endmodule
